module execute_tv();
endmodule