module fetch_tb();
endmodule